module top;

bit CLK = '0;
bit MNMX = '1;
bit TEST = '1;
bit RESET = '0;
bit READY = '1;
bit NMI = '0;
bit INTR = '0;
bit HOLD = '0;

wire logic [7:0] AD;
logic [19:8] A;
logic HLDA;
logic IOM;
logic WR;
logic RD;
logic SSO;
logic INTA;
logic ALE;
logic DTR;
logic DEN;


logic [19:0] Address;
wire [7:0]  Data;

Intel8088 P(CLK, MNMX, TEST, RESET, READY, NMI, INTR, HOLD, AD, A, HLDA, IOM, WR, RD, SSO, INTA, ALE, DTR, DEN);
//fsm f(.CLK(CLK),.ALE(ALE),.RD(RD),.WR(WR),.Address(Address),.RESET(RESET),.Data(Data));
//memory_2421 m(.Data(Data));
memory_1 m1(.CLK(CLK),.ALE(ALE),.IOM(IOM),.RD(RD),.WR(WR),.Data(Data),.Address(Address),.RESET(RESET));
memory_2 m2(.CLK(CLK),.ALE(ALE),.IOM(IOM),.RD(RD),.WR(WR),.Data(Data),.Address(Address),.RESET(RESET));
io_1 i1(.CLK(CLK),.ALE(ALE),.IOM(IOM),.RD(RD),.WR(WR),.Data(Data),.Address(Address),.RESET(RESET));
io_2 i2(.CLK(CLK),.ALE(ALE),.IOM(IOM),.RD(RD),.WR(WR),.Data(Data),.Address(Address),.RESET(RESET));
// 8282 Latch to latch bus address
always_latch
begin
if (ALE)
	Address <= {A, AD};
end

// 8286 transceiver
assign Data =  (DTR & ~DEN) ? AD   : 'z;
assign AD   = (~DTR & ~DEN) ? Data : 'z;


always #50 CLK = ~CLK;

initial
begin
$dumpfile("dump.vcd"); $dumpvars;

repeat (2) @(posedge CLK);
RESET = '1;
repeat (5) @(posedge CLK);
RESET = '0;

repeat(10000) @(posedge CLK);
$finish();
end

endmodule
